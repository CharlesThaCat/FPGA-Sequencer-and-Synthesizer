----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2018/06/11 17:59:10
-- Design Name: 
-- Module Name: sine_wave - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity sine_wave is
    Port ( clk_sw : in STD_LOGIC;
           dataout : out STD_LOGIC_VECTOR (7 downto 0));
end sine_wave;

architecture Behavioral of sine_wave is

signal index, index_next : integer range 0 to 628 := 0;
type memory_type is array (0 to 628) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
signal sine : memory_type := (128,129,131,132,133,134,136,137,138,140,141,142,143,145,146,147,148,150,151,152,153,155,156,157,158,160,161,162,163,165,166,167,168,169,171,172,173,174,175,177,178,179,180,181,183,184,185,186,187,188,189,190,192,193,194,195,196,197,198,199,200,201,202,203,204,205,206,207,208,209,210,211,212,213,214,215,216,217,218,219,220,221,222,222,223,224,225,226,227,227,228,229,230,231,231,232,233,234,234,235,236,236,237,238,238,239,240,240,241,241,242,243,243,244,244,245,245,246,246,247,247,248,248,249,249,249,250,250,251,251,251,252,252,252,253,253,253,253,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,255,254,254,254,254,253,253,253,253,252,252,252,251,251,251,250,250,250,249,249,248,248,247,247,246,246,245,245,244,244,243,243,242,242,241,240,240,239,238,238,237,237,236,235,234,234,233,232,231,231,230,229,228,228,227,226,225,224,223,223,222,221,220,219,218,217,216,215,214,214,213,212,211,210,209,208,207,206,205,204,203,201,200,199,198,197,196,195,194,193,192,191,190,188,187,186,185,184,183,182,180,179,178,177,176,174,173,172,171,170,168,167,166,165,164,162,161,160,159,157,156,155,154,152,151,150,149,147,146,145,144,142,141,140,138,137,136,135,133,132,131,129,128,127,126,124,123,122,121,119,118,117,115,114,113,112,110,109,108,107,105,104,103,102,100,99,98,97,95,94,93,92,90,89,88,87,86,84,83,82,81,80,78,77,76,75,74,73,71,70,69,68,67,66,65,63,62,61,60,59,58,57,56,55,54,53,52,51,50,49,48,47,46,45,44,43,42,41,40,39,38,37,36,35,35,34,33,32,31,30,29,29,28,27,26,26,25,24,23,23,22,21,20,20,19,18,18,17,16,16,15,15,14,13,13,12,12,11,11,10,10,9,9,8,8,7,7,7,6,6,5,5,5,4,4,4,3,3,3,3,2,2,2,2,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,2,2,2,2,2,3,3,3,4,4,4,5,5,5,6,6,6,7,7,8,8,9,9,9,10,10,11,12,12,13,13,14,14,15,16,16,17,17,18,19,19,20,21,21,22,23,24,24,25,26,27,27,28,29,30,31,32,32,33,34,35,36,37,38,39,40,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,58,59,60,61,62,63,64,65,66,67,69,70,71,72,73,74,75,77,78,79,80,81,83,84,85,86,87,89,90,91,92,93,95,96,97,98,100,101,102,103,105,106,107,108,110,111,112,114,115,116,117,119,120,121,122,124,125,126,128);


begin

process(clk_sw)
begin
  --to check the rising edge of the clock signal
if(rising_edge(clk_sw)) then     
    dataout <= std_logic_vector(to_unsigned(sine(index),8));
    index <= index_next;
end if;
end process;

index_next <= 0 when index = 628 else index + 1;


end Behavioral;
