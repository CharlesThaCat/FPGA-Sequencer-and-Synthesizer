----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2018/06/11 17:59:10
-- Design Name: 
-- Module Name: sine_wave - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity sine_wave is
    Port ( clk_sw_in : in STD_LOGIC;
           tone : in std_logic_vector (3 downto 0);
           clk_div_out : out STD_LOGIC;
           dataout : out STD_LOGIC_VECTOR (7 downto 0));
end sine_wave;

architecture Behavioral of sine_wave is

signal counter_phys_max : integer := 51;
signal clk_sw, clk_sw_tmp : STD_LOGIC := '0';

signal index, index_next, max_index: integer range 0 to 511 := 0;
signal counter_div, counter_div_next, counter_div_max: integer range 1 to 8 := 2;
signal clk_div: STD_LOGIC := '0';
type memory_type is array (0 to 511) of integer range 0 to 255; 
--ROM for storing the sine values generated by MATLAB.
signal A : memory_type := (127,130,132,135,138,140,143,145,148,151,153,156,158,161,164,166,169,171,174,176,178,181,183,186,188,190,193,195,197,199,201,204,206,208,210,212,214,216,218,219,221,223,225,226,228,230,231,233,234,236,237,238,240,241,242,243,244,245,246,247,248,249,250,250,251,252,252,253,253,254,254,254,255,255,255,255,255,255,255,255,255,254,254,254,253,253,252,252,251,250,250,249,248,247,246,245,244,243,242,241,240,238,237,236,234,233,231,230,228,226,225,223,221,219,217,216,214,212,210,208,205,203,201,199,197,195,192,190,188,185,183,181,178,176,173,171,168,166,163,161,158,156,153,150,148,145,143,140,137,135,132,129,127,124,121,119,116,114,111,108,106,103,101,98,95,93,90,88,85,83,80,78,75,73,71,68,66,64,61,59,57,55,52,50,48,46,44,42,40,38,36,34,33,31,29,27,26,24,23,21,20,18,17,16,14,13,12,11,10,9,8,7,6,5,4,4,3,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,2,3,4,4,5,6,7,8,9,10,11,12,13,15,16,17,19,20,22,23,25,26,28,30,31,33,35,37,39,41,43,45,47,49,51,53,55,57,60,62,64,66,69,71,74,76,78,81,83,86,88,91,93,96,99,101,104,106,109,112,114,117,119,122,125,127,130,133,135,138,141,143,146,148,151,154,156,159,161,164,166,169,171,174,176,179,181,184,186,188,191,193,195,197,200,202,204,206,208,210,212,214,216,218,220,221,223,225,227,228,230,231,233,234,236,237,239,240,241,242,243,244,245,246,247,248,249,250,251,251,252,252,253,253,254,254,254,255,255,255,255,255,255,255,255,255,254,254,254,253,253,252,252,251,250,250,249,248,247,246,245,244,243,242,241,239,238,237,235,234,232,231,229,228,226,224,223,221,219,217,215,213,211,209,207,205,203,201,199,197,194,192,190,187,185,183,180,178,175,173,170,168,165,163,160,158,155,153,150,147,145,142,140,137,134,132,129,126,124,121,118,116,113,111,108,105,103,100,98,95,92,90,87,85,82,80,77,75,73,70,68,65,63,61,59,56,54,52,50,48,46,44,42,40,38,36,34,32,31,29,27,26,24,22,21,19,18,17,15,14,13,12,11);
signal G : memory_type := (127,129,132,134,136,139,141,143,146,148,150,153,155,157,160,162,164,166,169,171,173,175,177,180,182,184,186,188,190,192,194,196,198,200,202,204,206,208,209,211,213,215,216,218,220,221,223,224,226,227,229,230,232,233,234,236,237,238,239,240,241,242,243,244,245,246,247,248,249,249,250,251,251,252,252,253,253,254,254,254,254,255,255,255,255,255,255,255,255,255,255,254,254,254,253,253,253,252,251,251,250,250,249,248,247,247,246,245,244,243,242,241,240,239,237,236,235,234,232,231,230,228,227,225,224,222,221,219,217,216,214,212,210,209,207,205,203,201,199,197,195,193,191,189,187,185,183,181,179,176,174,172,170,168,165,163,161,159,156,154,152,149,147,145,142,140,138,135,133,131,128,126,124,121,119,116,114,112,109,107,105,102,100,98,96,93,91,89,87,84,82,80,78,76,73,71,69,67,65,63,61,59,57,55,53,51,49,47,45,44,42,40,38,37,35,33,32,30,29,27,26,24,23,22,20,19,18,17,15,14,13,12,11,10,9,8,7,7,6,5,4,4,3,3,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,2,3,3,4,5,5,6,7,8,9,10,11,12,13,14,15,16,17,18,20,21,22,24,25,26,28,29,31,33,34,36,37,39,41,43,44,46,48,50,52,54,56,58,60,62,64,66,68,70,72,74,76,79,81,83,85,87,90,92,94,97,99,101,103,106,108,110,113,115,117,120,122,125,127,129,132,134,136,139,141,143,146,148,150,153,155,157,160,162,164,166,169,171,173,175,177,180,182,184,186,188,190,192,194,196,198,200,202,204,206,208,209,211,213,215,216,218,220,221,223,224,226,227,229,230,232,233,234,236,237,238,239,240,241,242,243,244,245,246,247,248,249,249,250,251,251,252,252,253,253,254,254,254,254,255,255,255,255,255,255,255,255,255,255,254,254,254,253,253,253,252,252,251,250,250,249,248,247,247,246,245,244,243,242,241,240,239,238,236,235,234,232,231,230,228,227,225,224,222,221,219,217,216,214,212,211,209,207,205,203,201,199,197,195,193,191,189,187,185,183,181,179,177,174,172,170,168,165,163,161,159,156,154,152,149,147,145,142,140,138,135,133,131,128);
signal E : memory_type := (127,129,131,133,135,137,139,141,143,145,147,149,151,153,155,156,158,160,162,164,166,168,170,172,174,175,177,179,181,183,184,186,188,190,191,193,195,196,198,200,201,203,205,206,208,209,211,212,214,215,217,218,219,221,222,223,225,226,227,228,230,231,232,233,234,235,236,237,238,239,240,241,242,243,244,244,245,246,247,247,248,249,249,250,250,251,251,252,252,253,253,253,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,254,254,254,254,253,253,253,252,252,251,251,250,250,249,249,248,247,247,246,245,244,243,243,242,241,240,239,238,237,236,235,234,233,232,230,229,228,227,226,224,223,222,220,219,218,216,215,213,212,210,209,207,206,204,203,201,199,198,196,194,193,191,189,188,186,184,182,180,179,177,175,173,171,169,168,166,164,162,160,158,156,154,152,150,148,146,144,142,140,138,136,135,133,131,129,127,125,123,121,119,117,115,113,111,109,107,105,103,101,99,97,95,93,91,89,88,86,84,82,80,78,76,75,73,71,69,67,66,64,62,61,59,57,56,54,52,51,49,48,46,45,43,42,40,39,37,36,34,33,32,30,29,28,27,25,24,23,22,21,20,19,18,17,16,15,14,13,12,11,10,9,9,8,7,6,6,5,5,4,4,3,3,2,2,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,2,2,3,3,4,4,5,6,6,7,8,8,9,10,11,12,12,13,14,15,16,17,18,19,20,21,23,24,25,26,27,29,30,31,33,34,35,37,38,40,41,42,44,45,47,49,50,52,53,55,57,58,60,62,63,65,67,69,70,72,74,76,78,79,81,83,85,87,89,91,93,94,96,98,100,102,104,106,108,110,112,114,116,118,120,122,124,126,128,130,132,134,136,138,140,142,144,146,148,150,151,153,155,157,159,161,163,165,167,169,171,172,174,176,178,180,182,183,185,187,189,190,192,194,195,197,199,200,202,204,205,207,208,210,211,213,214,216,217,219,220,221,223,224,225,226,228,229,230,231,232,233,235,236,237,238,239,240,241,241,242,243,244,245,246,246,247,248,248,249,250,250,251,251,252,252,252,253,253,253,254,254,254,254,255,255,255,255,255,255,255,255,255,255);
signal D : memory_type := (127,129,131,132,134,136,138,139,141,143,145,146,148,150,152,153,155,157,158,160,162,164,165,167,169,170,172,174,175,177,178,180,182,183,185,186,188,190,191,193,194,196,197,199,200,201,203,204,206,207,208,210,211,213,214,215,216,218,219,220,221,222,224,225,226,227,228,229,230,231,232,233,234,235,236,237,238,239,240,241,241,242,243,244,244,245,246,246,247,248,248,249,249,250,250,251,251,252,252,252,253,253,253,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,254,254,254,254,253,253,253,253,252,252,251,251,251,250,250,249,249,248,247,247,246,245,245,244,243,243,242,241,240,239,239,238,237,236,235,234,233,232,231,230,229,228,227,226,224,223,222,221,220,218,217,216,215,213,212,211,209,208,207,205,204,202,201,199,198,197,195,194,192,191,189,187,186,184,183,181,180,178,176,175,173,171,170,168,166,165,163,161,160,158,156,154,153,151,149,147,146,144,142,140,139,137,135,133,132,130,128,126,125,123,121,119,118,116,114,112,110,109,107,105,104,102,100,98,97,95,93,91,90,88,86,85,83,81,80,78,77,75,73,72,70,69,67,65,64,62,61,59,58,56,55,53,52,51,49,48,46,45,44,42,41,40,38,37,36,35,33,32,31,30,29,28,27,25,24,23,22,21,20,19,18,17,17,16,15,14,13,12,12,11,10,9,9,8,7,7,6,6,5,5,4,4,3,3,2,2,2,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,8,8,9,10,10,11,12,12,13,14,15,16,17,18,19,19,20,21,22,23,25,26,27,28,29,30,31,32,34,35,36,37,39,40,41,42,44,45,47,48,49,51,52,54,55,57,58,59,61,63,64,66,67,69,70,72,73,75,77,78,80,82,83,85,87,88,90,92,93,95,97,99,100,102,104,105,107,109,111,112,114,116,118,119,121,123,125,127,128,130,132,134,135,137,139,141,142,144,146,148,149,151,153,155,156,158,160,161,163,165,167,168,170,172,173,175,176,178,180,181,183,184,186,188,189,191,192,194,195,197,198,200,201,203,204,205,207,208,210,211,212,213,215,216);
signal C : memory_type := (127,129,130,132,133,135,136,138,140,141,143,144,146,147,149,150,152,154,155,157,158,160,161,163,164,166,167,169,170,172,173,175,176,178,179,180,182,183,185,186,187,189,190,192,193,194,196,197,198,200,201,202,203,205,206,207,208,210,211,212,213,214,215,217,218,219,220,221,222,223,224,225,226,227,228,229,230,231,232,233,234,234,235,236,237,238,239,239,240,241,241,242,243,243,244,245,245,246,247,247,248,248,249,249,250,250,250,251,251,252,252,252,253,253,253,253,254,254,254,254,254,255,255,255,255,255,255,255,255,255,255,255,255,255,255,254,254,254,254,254,254,253,253,253,252,252,252,251,251,251,250,250,249,249,248,248,247,247,246,246,245,244,244,243,242,242,241,240,240,239,238,237,237,236,235,234,233,232,231,230,229,229,228,227,226,225,224,223,221,220,219,218,217,216,215,214,213,211,210,209,208,206,205,204,203,201,200,199,198,196,195,194,192,191,190,188,187,185,184,183,181,180,178,177,175,174,172,171,169,168,166,165,163,162,160,159,157,156,154,153,151,150,148,147,145,143,142,140,139,137,136,134,133,131,129,128,126,125,123,121,120,118,117,115,114,112,111,109,107,106,104,103,101,100,98,97,95,94,92,91,89,88,86,85,83,82,80,79,77,76,74,73,71,70,69,67,66,64,63,62,60,59,58,56,55,54,53,51,50,49,48,46,45,44,43,41,40,39,38,37,36,35,34,33,31,30,29,28,27,26,25,25,24,23,22,21,20,19,18,17,17,16,15,14,14,13,12,12,11,10,10,9,8,8,7,7,6,6,5,5,4,4,3,3,3,2,2,2,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,7,8,9,9,10,11,11,12,13,13,14,15,15,16,17,18,19,20,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,39,40,41,42,43,44,46,47,48,49,51,52,53,54,56,57,58,60,61,62,64,65,67,68,69,71,72,74,75,76,78,79,81,82,84,85,87,88,90,91,93,94,96,97,99,100,102,104,105,107,108,110,111,113,114,116,118,119,121,122,124,125,127);
signal wave : memory_type;
begin

-- divide input 100M clk, to fit the output physical frequency
my_div: process (clk_sw_in,clk_sw_tmp)              
variable div_cnt : integer := 0;   
 begin
    if (rising_edge(clk_sw_in)) then   
       if (div_cnt = counter_phys_max) then 
          clk_sw_tmp <= not clk_sw_tmp; 
          div_cnt := 0; 
       else
          div_cnt := div_cnt + 1; 
       end if; 
    end if; 
    clk_sw <= clk_sw_tmp; 
 end process my_div; 

-- predefine waveform values according to input tone pitch
process(clk_sw, tone)
begin
    case tone is
        when "0000" =>
            max_index <= 0;
            wave <= C;
        when "0001" => -- C4
            max_index <= 511;
            counter_div_max <= 8;
            wave <= C;
        when "0110" => -- C5
            max_index <= 511;
            counter_div_max <= 4;
            wave <= C;
        when "1011" => -- C6 
            max_index <= 511;
            wave <= C;
        when "0010" => -- D4
            max_index <= 455;
            counter_div_max <= 8;
            wave <= D;
        when "0111" => -- D5
            max_index <= 455;
            counter_div_max <= 4;
            wave <= D;
        when "1100" => -- D6 
            max_index <= 455;
            wave <= D;
        when "0011" => -- E4
            max_index <= 407;
            counter_div_max <= 8;
            wave <= E;
        when "1000" => -- E5
            max_index <= 407;
            counter_div_max <= 4;
            wave <= E;
        when "1101" => -- E6 
            max_index <= 407;
            wave <= E;
        when "0100" => -- G4
            max_index <= 342;
            counter_div_max <= 8;
            wave <= G;
        when "1001" => -- G5
            max_index <= 342;
            counter_div_max <= 4;
            wave <= G;
        when "1110" => -- G6 
            max_index <= 342;
            wave <= G;
        when "0101" => -- A4
            max_index <= 305;
            counter_div_max <= 8;
            wave <= A;
        when "1010" => -- A5
            max_index <= 305;
            counter_div_max <= 4;
            wave <= A;
        when "1111" => -- A6 
            max_index <= 305;
            wave <= A;
        when others =>
    end case;
end process;

-- frequency divider for octaves
process (clk_sw, counter_div_max)
begin
if (rising_edge(clk_sw)) then
    counter_div <= counter_div_next;
    if counter_div = 1 then
        clk_div <= '1';
    else
        clk_div <= '0';
    end if;
end if;
end process;
counter_div_next <= counter_div + 1 when counter_div < counter_div_max + 1 else 1;  

-- output value loader, reads the array waveform value 
process(clk_div)
begin
if(rising_edge(clk_div)) then     
    dataout <= std_logic_vector(to_unsigned(wave(index),8));
    index <= index_next;
end if;
end process;
index_next <= 0 when index = max_index else index + 1;

clk_div_out <= clk_div;
end Behavioral;
